library ieee;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

use IEEE.std_logic_arith.all;

entity LUT_MAC is
	PORT(  
	T:  IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	Y:	IN STD_LOGIC_VECTOR(35 DOWNTO 0);
	I:	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	X:	OUT STD_LOGIC_VECTOR(35 DOWNTO 0);
	COEF:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
end LUT_MAC;

architecture LUT_MAC of LUT_MAC is	  
--COEFICIENTES
SIGNAL A0: STD_LOGIC_VECTOR(35 DOWNTO 0):="000000000000000000001100100110011000";
SIGNAL A1: STD_LOGIC_VECTOR(35 DOWNTO 0):="111111111111111110000011100000110101";
SIGNAL A2: STD_LOGIC_VECTOR(35 DOWNTO 0):="111111111111100001000000000110000010";
SIGNAL A3: STD_LOGIC_VECTOR(35 DOWNTO 0):="000000001000010101110110110011001110";
SIGNAL A4: STD_LOGIC_VECTOR(35 DOWNTO 0):="111111011011100101100010100011001100";
SIGNAL A5: STD_LOGIC_VECTOR(35 DOWNTO 0):="111111101101001100111000111101111010";
SIGNAL A6: STD_LOGIC_VECTOR(35 DOWNTO 0):="000111111111100101110010010001110100";
SIGNAL A7: STD_LOGIC_VECTOR(35 DOWNTO 0):="010000000101100001111001001111011110";

begin
	PROCESS(I)
	BEGIN
		CASE I IS
			WHEN "0000"=>	--0
			   X<=A0;	
			COEF<=T;
			WHEN "0001"=>	--1
			   X<=A1;
			COEF<="00010000";	--1
			WHEN "0010"=>	--0
			   X<=Y;
			COEF<=T;
			WHEN "0011"=>	--1
			   X<=A2;
			COEF<="00010000";	--1
			WHEN "0100"=>	--0
			   X<=Y;
			COEF<=T;
			WHEN "0101"=>	--1
			   X<=A3;
			COEF<="00010000";	--1
			WHEN "0110"=>	--0
			   X<=Y;
			COEF<=T;
			WHEN "0111"=>	--1
			   X<=A4;
			COEF<="00010000";	--1
			WHEN "1000"=>	--0
			   X<=Y;
			COEF<=T;
			WHEN "1001"=>	--1
			   X<=A5;
			COEF<="00010000";	--1
			WHEN "1010"=>	--0
			   X<=Y;
			COEF<=T;
			WHEN "1011"=>	--1
			   X<=A6;
			COEF<="00010000";	--1
			WHEN "1100"=>	--0
			   X<=Y;
			COEF<=T;
			WHEN "1101"=>	--1
			   X<=A7;
			COEF<="00010000";	--1		  
			WHEN OTHERS=>
			   X<=A0;	
			COEF<=T;
		END CASE;
	END PROCESS;
end LUT_MAC;
